module twoscompliment(
    input A0, A1, A2, A3, B0, B1, B2, B3, 
   
    output Twos0, Twos1, Twos2, Twos3, Twos4, Twos5, Twos6, Twos7 
);






endmodule